
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hd87ba53f;
    ram_cell[       1] = 32'h0;  // 32'ha7e94b71;
    ram_cell[       2] = 32'h0;  // 32'hdca627fd;
    ram_cell[       3] = 32'h0;  // 32'h04b27f41;
    ram_cell[       4] = 32'h0;  // 32'h2fa7318e;
    ram_cell[       5] = 32'h0;  // 32'hecda1d9d;
    ram_cell[       6] = 32'h0;  // 32'he4289508;
    ram_cell[       7] = 32'h0;  // 32'h6e1a59ce;
    ram_cell[       8] = 32'h0;  // 32'hc967e790;
    ram_cell[       9] = 32'h0;  // 32'h8be278c6;
    ram_cell[      10] = 32'h0;  // 32'hbef65710;
    ram_cell[      11] = 32'h0;  // 32'hcf778b95;
    ram_cell[      12] = 32'h0;  // 32'h63836ddf;
    ram_cell[      13] = 32'h0;  // 32'h0be78b01;
    ram_cell[      14] = 32'h0;  // 32'h2aa249d1;
    ram_cell[      15] = 32'h0;  // 32'h30c46603;
    ram_cell[      16] = 32'h0;  // 32'h79a6e41c;
    ram_cell[      17] = 32'h0;  // 32'h7ba60e3d;
    ram_cell[      18] = 32'h0;  // 32'hcf73d53d;
    ram_cell[      19] = 32'h0;  // 32'h3a55e73c;
    ram_cell[      20] = 32'h0;  // 32'h0d9eeac9;
    ram_cell[      21] = 32'h0;  // 32'ha71e4bd9;
    ram_cell[      22] = 32'h0;  // 32'h411c3471;
    ram_cell[      23] = 32'h0;  // 32'hec135fa4;
    ram_cell[      24] = 32'h0;  // 32'h68eba929;
    ram_cell[      25] = 32'h0;  // 32'hbe9427f7;
    ram_cell[      26] = 32'h0;  // 32'h09827d08;
    ram_cell[      27] = 32'h0;  // 32'hff1feed7;
    ram_cell[      28] = 32'h0;  // 32'h73f799e8;
    ram_cell[      29] = 32'h0;  // 32'h775b9b89;
    ram_cell[      30] = 32'h0;  // 32'hb6806d35;
    ram_cell[      31] = 32'h0;  // 32'hf08b7a5f;
    ram_cell[      32] = 32'h0;  // 32'h6ce3b804;
    ram_cell[      33] = 32'h0;  // 32'hf48d9c44;
    ram_cell[      34] = 32'h0;  // 32'hee36ed46;
    ram_cell[      35] = 32'h0;  // 32'hd672d722;
    ram_cell[      36] = 32'h0;  // 32'h75b30564;
    ram_cell[      37] = 32'h0;  // 32'h02209760;
    ram_cell[      38] = 32'h0;  // 32'hc17d4f61;
    ram_cell[      39] = 32'h0;  // 32'h7d1bdff2;
    ram_cell[      40] = 32'h0;  // 32'he09c9adf;
    ram_cell[      41] = 32'h0;  // 32'h84a3c846;
    ram_cell[      42] = 32'h0;  // 32'hd154010c;
    ram_cell[      43] = 32'h0;  // 32'h95309926;
    ram_cell[      44] = 32'h0;  // 32'h0e14f8e2;
    ram_cell[      45] = 32'h0;  // 32'he3463ff8;
    ram_cell[      46] = 32'h0;  // 32'hd3eff2e8;
    ram_cell[      47] = 32'h0;  // 32'h12f89b13;
    ram_cell[      48] = 32'h0;  // 32'hcaf88031;
    ram_cell[      49] = 32'h0;  // 32'hbb85b2d2;
    ram_cell[      50] = 32'h0;  // 32'h28ff45f0;
    ram_cell[      51] = 32'h0;  // 32'h9c216cf6;
    ram_cell[      52] = 32'h0;  // 32'h70a91430;
    ram_cell[      53] = 32'h0;  // 32'h99a11abf;
    ram_cell[      54] = 32'h0;  // 32'he904f01c;
    ram_cell[      55] = 32'h0;  // 32'he95b4d57;
    ram_cell[      56] = 32'h0;  // 32'h20195106;
    ram_cell[      57] = 32'h0;  // 32'h1da2877f;
    ram_cell[      58] = 32'h0;  // 32'h17994a53;
    ram_cell[      59] = 32'h0;  // 32'he47fb07a;
    ram_cell[      60] = 32'h0;  // 32'h6db45f0d;
    ram_cell[      61] = 32'h0;  // 32'h076f3e98;
    ram_cell[      62] = 32'h0;  // 32'hf867d99b;
    ram_cell[      63] = 32'h0;  // 32'h91245070;
    ram_cell[      64] = 32'h0;  // 32'hb290a532;
    ram_cell[      65] = 32'h0;  // 32'hbc0b0364;
    ram_cell[      66] = 32'h0;  // 32'h956eb258;
    ram_cell[      67] = 32'h0;  // 32'h45944b3c;
    ram_cell[      68] = 32'h0;  // 32'h06bc0b50;
    ram_cell[      69] = 32'h0;  // 32'h0dc2f594;
    ram_cell[      70] = 32'h0;  // 32'h13c576ef;
    ram_cell[      71] = 32'h0;  // 32'ha7b288ac;
    ram_cell[      72] = 32'h0;  // 32'hc30bc738;
    ram_cell[      73] = 32'h0;  // 32'h79eba97d;
    ram_cell[      74] = 32'h0;  // 32'h3fe90a74;
    ram_cell[      75] = 32'h0;  // 32'h952d3d2b;
    ram_cell[      76] = 32'h0;  // 32'h0efaf073;
    ram_cell[      77] = 32'h0;  // 32'hbdb6bc0a;
    ram_cell[      78] = 32'h0;  // 32'h26702e5f;
    ram_cell[      79] = 32'h0;  // 32'h14a64e95;
    ram_cell[      80] = 32'h0;  // 32'h3a28aa6e;
    ram_cell[      81] = 32'h0;  // 32'hbf716301;
    ram_cell[      82] = 32'h0;  // 32'h05dbd5f2;
    ram_cell[      83] = 32'h0;  // 32'h36e5697e;
    ram_cell[      84] = 32'h0;  // 32'hcf2df09c;
    ram_cell[      85] = 32'h0;  // 32'hf2d58bde;
    ram_cell[      86] = 32'h0;  // 32'hc13a2cf0;
    ram_cell[      87] = 32'h0;  // 32'h2fde4f8c;
    ram_cell[      88] = 32'h0;  // 32'h4235af04;
    ram_cell[      89] = 32'h0;  // 32'h0edbd476;
    ram_cell[      90] = 32'h0;  // 32'h9dee35e1;
    ram_cell[      91] = 32'h0;  // 32'he75e14ff;
    ram_cell[      92] = 32'h0;  // 32'h9a61485a;
    ram_cell[      93] = 32'h0;  // 32'h7cfb2ca5;
    ram_cell[      94] = 32'h0;  // 32'h392b7bd1;
    ram_cell[      95] = 32'h0;  // 32'h70ab2efa;
    ram_cell[      96] = 32'h0;  // 32'hd903bae9;
    ram_cell[      97] = 32'h0;  // 32'h8b508610;
    ram_cell[      98] = 32'h0;  // 32'hbb5822fe;
    ram_cell[      99] = 32'h0;  // 32'hb2e4421f;
    ram_cell[     100] = 32'h0;  // 32'h56e3f59d;
    ram_cell[     101] = 32'h0;  // 32'hab5fa394;
    ram_cell[     102] = 32'h0;  // 32'hf7e05cc7;
    ram_cell[     103] = 32'h0;  // 32'hf10eadb9;
    ram_cell[     104] = 32'h0;  // 32'h92fdc1a2;
    ram_cell[     105] = 32'h0;  // 32'h05d7238d;
    ram_cell[     106] = 32'h0;  // 32'h1575c568;
    ram_cell[     107] = 32'h0;  // 32'h32f1fdb6;
    ram_cell[     108] = 32'h0;  // 32'h3328e100;
    ram_cell[     109] = 32'h0;  // 32'h99979dfd;
    ram_cell[     110] = 32'h0;  // 32'h6f4fbb8b;
    ram_cell[     111] = 32'h0;  // 32'h68c6c116;
    ram_cell[     112] = 32'h0;  // 32'ha08d57f1;
    ram_cell[     113] = 32'h0;  // 32'he20df008;
    ram_cell[     114] = 32'h0;  // 32'h28124e59;
    ram_cell[     115] = 32'h0;  // 32'h6d0a052b;
    ram_cell[     116] = 32'h0;  // 32'hd56b0572;
    ram_cell[     117] = 32'h0;  // 32'h0f5e53d2;
    ram_cell[     118] = 32'h0;  // 32'hb7bbffa9;
    ram_cell[     119] = 32'h0;  // 32'h3bad1b24;
    ram_cell[     120] = 32'h0;  // 32'h25bb1726;
    ram_cell[     121] = 32'h0;  // 32'h272fcc52;
    ram_cell[     122] = 32'h0;  // 32'hce7c7b70;
    ram_cell[     123] = 32'h0;  // 32'hb5a7660f;
    ram_cell[     124] = 32'h0;  // 32'h88cce636;
    ram_cell[     125] = 32'h0;  // 32'h5d8f7a11;
    ram_cell[     126] = 32'h0;  // 32'hdc25119c;
    ram_cell[     127] = 32'h0;  // 32'h96e96719;
    ram_cell[     128] = 32'h0;  // 32'hd98beb5d;
    ram_cell[     129] = 32'h0;  // 32'h114f4dba;
    ram_cell[     130] = 32'h0;  // 32'hb511745d;
    ram_cell[     131] = 32'h0;  // 32'hdd95be40;
    ram_cell[     132] = 32'h0;  // 32'hda43b432;
    ram_cell[     133] = 32'h0;  // 32'h17afe10b;
    ram_cell[     134] = 32'h0;  // 32'hf145651a;
    ram_cell[     135] = 32'h0;  // 32'h8d34244d;
    ram_cell[     136] = 32'h0;  // 32'h80b866c7;
    ram_cell[     137] = 32'h0;  // 32'h13f0385e;
    ram_cell[     138] = 32'h0;  // 32'hc5853fd7;
    ram_cell[     139] = 32'h0;  // 32'hc6aa61cc;
    ram_cell[     140] = 32'h0;  // 32'he53d914d;
    ram_cell[     141] = 32'h0;  // 32'hca7c587b;
    ram_cell[     142] = 32'h0;  // 32'hb80fa06d;
    ram_cell[     143] = 32'h0;  // 32'hb415cfdf;
    ram_cell[     144] = 32'h0;  // 32'h31a28c8c;
    ram_cell[     145] = 32'h0;  // 32'hb5738f49;
    ram_cell[     146] = 32'h0;  // 32'h84057251;
    ram_cell[     147] = 32'h0;  // 32'h0536d2d1;
    ram_cell[     148] = 32'h0;  // 32'h099bebbd;
    ram_cell[     149] = 32'h0;  // 32'h089cffa5;
    ram_cell[     150] = 32'h0;  // 32'h113e7965;
    ram_cell[     151] = 32'h0;  // 32'h5a2355e1;
    ram_cell[     152] = 32'h0;  // 32'h60de37cb;
    ram_cell[     153] = 32'h0;  // 32'hc22aabe4;
    ram_cell[     154] = 32'h0;  // 32'h1115ef48;
    ram_cell[     155] = 32'h0;  // 32'h1ad79259;
    ram_cell[     156] = 32'h0;  // 32'h2f0b64b1;
    ram_cell[     157] = 32'h0;  // 32'h8903e171;
    ram_cell[     158] = 32'h0;  // 32'h4cf87834;
    ram_cell[     159] = 32'h0;  // 32'h757f48db;
    ram_cell[     160] = 32'h0;  // 32'h917d6a9f;
    ram_cell[     161] = 32'h0;  // 32'h892e3923;
    ram_cell[     162] = 32'h0;  // 32'h492a563f;
    ram_cell[     163] = 32'h0;  // 32'hfd3bef88;
    ram_cell[     164] = 32'h0;  // 32'h054c0511;
    ram_cell[     165] = 32'h0;  // 32'hdd2581b7;
    ram_cell[     166] = 32'h0;  // 32'h75040f3a;
    ram_cell[     167] = 32'h0;  // 32'h9c9f42c2;
    ram_cell[     168] = 32'h0;  // 32'h03493acf;
    ram_cell[     169] = 32'h0;  // 32'h8eac1331;
    ram_cell[     170] = 32'h0;  // 32'hbcc916bc;
    ram_cell[     171] = 32'h0;  // 32'hc50d3aa0;
    ram_cell[     172] = 32'h0;  // 32'h7eaceede;
    ram_cell[     173] = 32'h0;  // 32'h49f8d823;
    ram_cell[     174] = 32'h0;  // 32'h0cee355e;
    ram_cell[     175] = 32'h0;  // 32'h0218e3a7;
    ram_cell[     176] = 32'h0;  // 32'h19869183;
    ram_cell[     177] = 32'h0;  // 32'hb065887b;
    ram_cell[     178] = 32'h0;  // 32'he8441a3f;
    ram_cell[     179] = 32'h0;  // 32'h9ca94dfe;
    ram_cell[     180] = 32'h0;  // 32'h73745029;
    ram_cell[     181] = 32'h0;  // 32'h499ecf44;
    ram_cell[     182] = 32'h0;  // 32'he5601649;
    ram_cell[     183] = 32'h0;  // 32'hbb0ee942;
    ram_cell[     184] = 32'h0;  // 32'h48a6b48b;
    ram_cell[     185] = 32'h0;  // 32'hea3853e8;
    ram_cell[     186] = 32'h0;  // 32'h0de001cb;
    ram_cell[     187] = 32'h0;  // 32'h2a6e6af5;
    ram_cell[     188] = 32'h0;  // 32'hf8158201;
    ram_cell[     189] = 32'h0;  // 32'h5c6e5da2;
    ram_cell[     190] = 32'h0;  // 32'h5e1b2fcb;
    ram_cell[     191] = 32'h0;  // 32'hd8722353;
    ram_cell[     192] = 32'h0;  // 32'h502c96d9;
    ram_cell[     193] = 32'h0;  // 32'h17fc26c5;
    ram_cell[     194] = 32'h0;  // 32'h48293886;
    ram_cell[     195] = 32'h0;  // 32'h69de4988;
    ram_cell[     196] = 32'h0;  // 32'h0d592fea;
    ram_cell[     197] = 32'h0;  // 32'h20742a34;
    ram_cell[     198] = 32'h0;  // 32'h6debc8fe;
    ram_cell[     199] = 32'h0;  // 32'hdbbf4375;
    ram_cell[     200] = 32'h0;  // 32'hb0dd5adb;
    ram_cell[     201] = 32'h0;  // 32'hc1c833b3;
    ram_cell[     202] = 32'h0;  // 32'h6c96f671;
    ram_cell[     203] = 32'h0;  // 32'h952248db;
    ram_cell[     204] = 32'h0;  // 32'h51b2c3fc;
    ram_cell[     205] = 32'h0;  // 32'h6a9cd213;
    ram_cell[     206] = 32'h0;  // 32'h608b88aa;
    ram_cell[     207] = 32'h0;  // 32'h53a5dec9;
    ram_cell[     208] = 32'h0;  // 32'hb21ac961;
    ram_cell[     209] = 32'h0;  // 32'h0172ca9c;
    ram_cell[     210] = 32'h0;  // 32'h96f5e146;
    ram_cell[     211] = 32'h0;  // 32'hc7b76b20;
    ram_cell[     212] = 32'h0;  // 32'h826393e9;
    ram_cell[     213] = 32'h0;  // 32'hbdedc59a;
    ram_cell[     214] = 32'h0;  // 32'h048a4290;
    ram_cell[     215] = 32'h0;  // 32'hb9faee30;
    ram_cell[     216] = 32'h0;  // 32'h517458b7;
    ram_cell[     217] = 32'h0;  // 32'h57701209;
    ram_cell[     218] = 32'h0;  // 32'h715e03f9;
    ram_cell[     219] = 32'h0;  // 32'h1f1920c8;
    ram_cell[     220] = 32'h0;  // 32'h634cd075;
    ram_cell[     221] = 32'h0;  // 32'h17687b7c;
    ram_cell[     222] = 32'h0;  // 32'hc6aca0d5;
    ram_cell[     223] = 32'h0;  // 32'h5d70c18e;
    ram_cell[     224] = 32'h0;  // 32'h34f413be;
    ram_cell[     225] = 32'h0;  // 32'hf69772b9;
    ram_cell[     226] = 32'h0;  // 32'h482a30a1;
    ram_cell[     227] = 32'h0;  // 32'h2db65ddc;
    ram_cell[     228] = 32'h0;  // 32'h2499846a;
    ram_cell[     229] = 32'h0;  // 32'h1b8e8c38;
    ram_cell[     230] = 32'h0;  // 32'h404c6eae;
    ram_cell[     231] = 32'h0;  // 32'hefa674de;
    ram_cell[     232] = 32'h0;  // 32'hb1e0bcc6;
    ram_cell[     233] = 32'h0;  // 32'hfbd2cb24;
    ram_cell[     234] = 32'h0;  // 32'h79420844;
    ram_cell[     235] = 32'h0;  // 32'h3fd7b4ef;
    ram_cell[     236] = 32'h0;  // 32'h228317f1;
    ram_cell[     237] = 32'h0;  // 32'hfdcf1956;
    ram_cell[     238] = 32'h0;  // 32'h6321ca18;
    ram_cell[     239] = 32'h0;  // 32'h10486c98;
    ram_cell[     240] = 32'h0;  // 32'h4c16785e;
    ram_cell[     241] = 32'h0;  // 32'h47d715f9;
    ram_cell[     242] = 32'h0;  // 32'h4039cbb3;
    ram_cell[     243] = 32'h0;  // 32'h2f4a651f;
    ram_cell[     244] = 32'h0;  // 32'h40689750;
    ram_cell[     245] = 32'h0;  // 32'h6bee5c1b;
    ram_cell[     246] = 32'h0;  // 32'he756498c;
    ram_cell[     247] = 32'h0;  // 32'h56349b41;
    ram_cell[     248] = 32'h0;  // 32'h09f29156;
    ram_cell[     249] = 32'h0;  // 32'h67111ea5;
    ram_cell[     250] = 32'h0;  // 32'hbbb38c9d;
    ram_cell[     251] = 32'h0;  // 32'h29c7e4f3;
    ram_cell[     252] = 32'h0;  // 32'ha601d5cd;
    ram_cell[     253] = 32'h0;  // 32'hdedba696;
    ram_cell[     254] = 32'h0;  // 32'h65c079e0;
    ram_cell[     255] = 32'h0;  // 32'hd5961946;
    // src matrix A
    ram_cell[     256] = 32'hd90c1519;
    ram_cell[     257] = 32'hd578fbdd;
    ram_cell[     258] = 32'h07d68cc0;
    ram_cell[     259] = 32'h0efa386c;
    ram_cell[     260] = 32'h4e592452;
    ram_cell[     261] = 32'h52b45082;
    ram_cell[     262] = 32'hf7a2cb5d;
    ram_cell[     263] = 32'h27996286;
    ram_cell[     264] = 32'h2f36d4cd;
    ram_cell[     265] = 32'h67595722;
    ram_cell[     266] = 32'hee8b3841;
    ram_cell[     267] = 32'h68607a98;
    ram_cell[     268] = 32'h87059357;
    ram_cell[     269] = 32'hf1de4154;
    ram_cell[     270] = 32'hdc007aea;
    ram_cell[     271] = 32'h9f484ebb;
    ram_cell[     272] = 32'h766fe24b;
    ram_cell[     273] = 32'h4d9575e7;
    ram_cell[     274] = 32'h7979ce4b;
    ram_cell[     275] = 32'h18765000;
    ram_cell[     276] = 32'hfdc5b5c2;
    ram_cell[     277] = 32'hb917e186;
    ram_cell[     278] = 32'h47362d22;
    ram_cell[     279] = 32'h91db838f;
    ram_cell[     280] = 32'h7f58ee1a;
    ram_cell[     281] = 32'h4b2f8fc6;
    ram_cell[     282] = 32'he4cac9c0;
    ram_cell[     283] = 32'hd944fe24;
    ram_cell[     284] = 32'hda6fdaf7;
    ram_cell[     285] = 32'h3060ae51;
    ram_cell[     286] = 32'hd178a7c9;
    ram_cell[     287] = 32'h824fb258;
    ram_cell[     288] = 32'hce725642;
    ram_cell[     289] = 32'h09db5444;
    ram_cell[     290] = 32'h7f5f89c3;
    ram_cell[     291] = 32'h75439874;
    ram_cell[     292] = 32'hfed47313;
    ram_cell[     293] = 32'h346612fb;
    ram_cell[     294] = 32'hb3ccd152;
    ram_cell[     295] = 32'h3316e7a4;
    ram_cell[     296] = 32'hdbf92937;
    ram_cell[     297] = 32'h96f9a0c9;
    ram_cell[     298] = 32'h51ae05cf;
    ram_cell[     299] = 32'h8da363c2;
    ram_cell[     300] = 32'h466452f6;
    ram_cell[     301] = 32'h9fd41901;
    ram_cell[     302] = 32'hb2ed89dd;
    ram_cell[     303] = 32'hedb0199a;
    ram_cell[     304] = 32'h65c10e86;
    ram_cell[     305] = 32'h55e46c9d;
    ram_cell[     306] = 32'h5112b3c1;
    ram_cell[     307] = 32'hd0ce808a;
    ram_cell[     308] = 32'h038a5fee;
    ram_cell[     309] = 32'hffc1b65b;
    ram_cell[     310] = 32'h61555598;
    ram_cell[     311] = 32'h9641f202;
    ram_cell[     312] = 32'hb759ec9d;
    ram_cell[     313] = 32'h286dff7d;
    ram_cell[     314] = 32'hc1b18e7b;
    ram_cell[     315] = 32'hb46147d6;
    ram_cell[     316] = 32'ha28fc6ef;
    ram_cell[     317] = 32'h6f3f1f39;
    ram_cell[     318] = 32'hfa1f4546;
    ram_cell[     319] = 32'h9c649fce;
    ram_cell[     320] = 32'hdc405a1e;
    ram_cell[     321] = 32'hd0dcda09;
    ram_cell[     322] = 32'haa1b4218;
    ram_cell[     323] = 32'he4eee767;
    ram_cell[     324] = 32'hcc40b711;
    ram_cell[     325] = 32'hf15b7480;
    ram_cell[     326] = 32'h198c4480;
    ram_cell[     327] = 32'h11f44d53;
    ram_cell[     328] = 32'hbd705119;
    ram_cell[     329] = 32'hab7794fc;
    ram_cell[     330] = 32'h973d4415;
    ram_cell[     331] = 32'h7d806b29;
    ram_cell[     332] = 32'h1f44992e;
    ram_cell[     333] = 32'habcd066c;
    ram_cell[     334] = 32'h68be99a5;
    ram_cell[     335] = 32'hd0aec5f5;
    ram_cell[     336] = 32'h7d9bad60;
    ram_cell[     337] = 32'h7dc81376;
    ram_cell[     338] = 32'hc3a710d0;
    ram_cell[     339] = 32'he43bf95e;
    ram_cell[     340] = 32'h03726ad9;
    ram_cell[     341] = 32'h659d8022;
    ram_cell[     342] = 32'h857575d5;
    ram_cell[     343] = 32'h80f0aa09;
    ram_cell[     344] = 32'h4abc64f5;
    ram_cell[     345] = 32'hfbedb03f;
    ram_cell[     346] = 32'h8b697b60;
    ram_cell[     347] = 32'he77e35f7;
    ram_cell[     348] = 32'h76d3803f;
    ram_cell[     349] = 32'h693be00d;
    ram_cell[     350] = 32'h11435243;
    ram_cell[     351] = 32'hd290645e;
    ram_cell[     352] = 32'h2fa2c30d;
    ram_cell[     353] = 32'h4db52bca;
    ram_cell[     354] = 32'h7c27f2e1;
    ram_cell[     355] = 32'h04d264cf;
    ram_cell[     356] = 32'h184f1ec8;
    ram_cell[     357] = 32'hb86b10dd;
    ram_cell[     358] = 32'h48e08ead;
    ram_cell[     359] = 32'h89913178;
    ram_cell[     360] = 32'h9c21e7f7;
    ram_cell[     361] = 32'h6beff79a;
    ram_cell[     362] = 32'h04aede70;
    ram_cell[     363] = 32'hf73cc463;
    ram_cell[     364] = 32'hf2dc4f8f;
    ram_cell[     365] = 32'hc015a93e;
    ram_cell[     366] = 32'hc8b25840;
    ram_cell[     367] = 32'h8b6aed30;
    ram_cell[     368] = 32'he4782e27;
    ram_cell[     369] = 32'hc665bb4f;
    ram_cell[     370] = 32'h65b8065a;
    ram_cell[     371] = 32'hc6779651;
    ram_cell[     372] = 32'hea8fc9b6;
    ram_cell[     373] = 32'h1a17ea22;
    ram_cell[     374] = 32'h45aabbcb;
    ram_cell[     375] = 32'hc23b135d;
    ram_cell[     376] = 32'h51930076;
    ram_cell[     377] = 32'h431393c1;
    ram_cell[     378] = 32'hbf5e426e;
    ram_cell[     379] = 32'hf330ac7d;
    ram_cell[     380] = 32'hf1fcc2cd;
    ram_cell[     381] = 32'h9f2a0081;
    ram_cell[     382] = 32'h2082e7c5;
    ram_cell[     383] = 32'he2536bc9;
    ram_cell[     384] = 32'h5442fa2b;
    ram_cell[     385] = 32'h1c0c5ead;
    ram_cell[     386] = 32'h578f0cec;
    ram_cell[     387] = 32'ha0d4b7ed;
    ram_cell[     388] = 32'hfb35107e;
    ram_cell[     389] = 32'h23886dad;
    ram_cell[     390] = 32'h963ddec7;
    ram_cell[     391] = 32'hd940643c;
    ram_cell[     392] = 32'h2b56e3c2;
    ram_cell[     393] = 32'h3919fa42;
    ram_cell[     394] = 32'hddc6cf76;
    ram_cell[     395] = 32'h4b8f0cf3;
    ram_cell[     396] = 32'h4f0b76f0;
    ram_cell[     397] = 32'h2e2f5f29;
    ram_cell[     398] = 32'h997e25fd;
    ram_cell[     399] = 32'h4a9ed9f3;
    ram_cell[     400] = 32'h4410fe29;
    ram_cell[     401] = 32'ha889970f;
    ram_cell[     402] = 32'hbd9e7ad3;
    ram_cell[     403] = 32'ha40cfd05;
    ram_cell[     404] = 32'ha1637829;
    ram_cell[     405] = 32'h0d447abf;
    ram_cell[     406] = 32'hd6508155;
    ram_cell[     407] = 32'h4efab885;
    ram_cell[     408] = 32'h57fe6169;
    ram_cell[     409] = 32'h08c13f76;
    ram_cell[     410] = 32'hcff168ff;
    ram_cell[     411] = 32'h115917bb;
    ram_cell[     412] = 32'hc1ecaf14;
    ram_cell[     413] = 32'h19723bc1;
    ram_cell[     414] = 32'ha55c1b97;
    ram_cell[     415] = 32'h090eb324;
    ram_cell[     416] = 32'h6d04c794;
    ram_cell[     417] = 32'hd9dfc6c4;
    ram_cell[     418] = 32'hc79ce213;
    ram_cell[     419] = 32'h70a7f80d;
    ram_cell[     420] = 32'hbdeb6835;
    ram_cell[     421] = 32'h942dc9a8;
    ram_cell[     422] = 32'hbd02a3f3;
    ram_cell[     423] = 32'h77ee371c;
    ram_cell[     424] = 32'h97ceed7d;
    ram_cell[     425] = 32'h1bd664de;
    ram_cell[     426] = 32'h9058ce38;
    ram_cell[     427] = 32'h1b5150d2;
    ram_cell[     428] = 32'he27b1820;
    ram_cell[     429] = 32'he8d3132a;
    ram_cell[     430] = 32'he30f4f2f;
    ram_cell[     431] = 32'ha46ab418;
    ram_cell[     432] = 32'h46e357c4;
    ram_cell[     433] = 32'h8831a5f8;
    ram_cell[     434] = 32'ha914b07e;
    ram_cell[     435] = 32'hc331762a;
    ram_cell[     436] = 32'h2b5e290e;
    ram_cell[     437] = 32'h9fd97720;
    ram_cell[     438] = 32'h8eb118ed;
    ram_cell[     439] = 32'he2ed9fb6;
    ram_cell[     440] = 32'h08a83bae;
    ram_cell[     441] = 32'h746c95fd;
    ram_cell[     442] = 32'h8353c80d;
    ram_cell[     443] = 32'h14e0f4ee;
    ram_cell[     444] = 32'hcf1d2ca5;
    ram_cell[     445] = 32'h2d492098;
    ram_cell[     446] = 32'hc91e33f5;
    ram_cell[     447] = 32'h2e2d4d10;
    ram_cell[     448] = 32'hd2f888b4;
    ram_cell[     449] = 32'h5af28fc3;
    ram_cell[     450] = 32'h88b2d2ce;
    ram_cell[     451] = 32'h81dead36;
    ram_cell[     452] = 32'hff142d87;
    ram_cell[     453] = 32'h9ef429bf;
    ram_cell[     454] = 32'h920a89e3;
    ram_cell[     455] = 32'hcd74c145;
    ram_cell[     456] = 32'h7965351d;
    ram_cell[     457] = 32'h6c35a0e1;
    ram_cell[     458] = 32'h04d8be0a;
    ram_cell[     459] = 32'hed9af081;
    ram_cell[     460] = 32'hdfbf1e8c;
    ram_cell[     461] = 32'h00d89920;
    ram_cell[     462] = 32'h7b74ac01;
    ram_cell[     463] = 32'h578da41f;
    ram_cell[     464] = 32'h3719c8e7;
    ram_cell[     465] = 32'h2ed18dd6;
    ram_cell[     466] = 32'hf67e8b8d;
    ram_cell[     467] = 32'h38b1fdb6;
    ram_cell[     468] = 32'h994b8869;
    ram_cell[     469] = 32'hbfdfab29;
    ram_cell[     470] = 32'hf3b26e1f;
    ram_cell[     471] = 32'h734863ad;
    ram_cell[     472] = 32'h9d46e179;
    ram_cell[     473] = 32'h8aa24836;
    ram_cell[     474] = 32'h61cc9d36;
    ram_cell[     475] = 32'h4d3c3e3f;
    ram_cell[     476] = 32'hf0328c96;
    ram_cell[     477] = 32'h7c4386ab;
    ram_cell[     478] = 32'hcf04ac31;
    ram_cell[     479] = 32'hedfe03a1;
    ram_cell[     480] = 32'h7804a637;
    ram_cell[     481] = 32'h641d30e5;
    ram_cell[     482] = 32'h7c386002;
    ram_cell[     483] = 32'h7ad0b875;
    ram_cell[     484] = 32'h611f962a;
    ram_cell[     485] = 32'hb81560a8;
    ram_cell[     486] = 32'ha6e01d93;
    ram_cell[     487] = 32'h5584aa89;
    ram_cell[     488] = 32'h7a2a6fdd;
    ram_cell[     489] = 32'h8dcee6cb;
    ram_cell[     490] = 32'haabb8344;
    ram_cell[     491] = 32'h19296a82;
    ram_cell[     492] = 32'h68d6a9fb;
    ram_cell[     493] = 32'hc38355fb;
    ram_cell[     494] = 32'h62a0c915;
    ram_cell[     495] = 32'h86ae88a8;
    ram_cell[     496] = 32'hd9819b62;
    ram_cell[     497] = 32'hacb408ed;
    ram_cell[     498] = 32'h85245efa;
    ram_cell[     499] = 32'hccf8531e;
    ram_cell[     500] = 32'h790ea2ba;
    ram_cell[     501] = 32'h2dd61436;
    ram_cell[     502] = 32'hd9f92ac0;
    ram_cell[     503] = 32'h21566a32;
    ram_cell[     504] = 32'h1083735e;
    ram_cell[     505] = 32'hb45110be;
    ram_cell[     506] = 32'h1eeb4665;
    ram_cell[     507] = 32'h25ba5b2f;
    ram_cell[     508] = 32'h39c164cb;
    ram_cell[     509] = 32'h7fe01b04;
    ram_cell[     510] = 32'h4937bd20;
    ram_cell[     511] = 32'h8c529218;
    // src matrix B
    ram_cell[     512] = 32'h028eea9b;
    ram_cell[     513] = 32'h071ca459;
    ram_cell[     514] = 32'h358e4414;
    ram_cell[     515] = 32'hb5933f8d;
    ram_cell[     516] = 32'h53757ef4;
    ram_cell[     517] = 32'h5fdf121c;
    ram_cell[     518] = 32'hcbe13b46;
    ram_cell[     519] = 32'h61a1cffa;
    ram_cell[     520] = 32'h537c7721;
    ram_cell[     521] = 32'h1da7454b;
    ram_cell[     522] = 32'h138b8cd2;
    ram_cell[     523] = 32'h98812a82;
    ram_cell[     524] = 32'h68111b60;
    ram_cell[     525] = 32'h06d3687a;
    ram_cell[     526] = 32'h82dd6bc1;
    ram_cell[     527] = 32'hd9afd7cb;
    ram_cell[     528] = 32'ha612ffb0;
    ram_cell[     529] = 32'h26e8fa4f;
    ram_cell[     530] = 32'h52036389;
    ram_cell[     531] = 32'h6aa26ffb;
    ram_cell[     532] = 32'ha2e6e995;
    ram_cell[     533] = 32'h3b9936c1;
    ram_cell[     534] = 32'hf0882721;
    ram_cell[     535] = 32'hcabdf86a;
    ram_cell[     536] = 32'h53739c5b;
    ram_cell[     537] = 32'h27ed641a;
    ram_cell[     538] = 32'hf0132caf;
    ram_cell[     539] = 32'h9294cedb;
    ram_cell[     540] = 32'h5fbdcfef;
    ram_cell[     541] = 32'h160531f2;
    ram_cell[     542] = 32'h760b7668;
    ram_cell[     543] = 32'h6d6e3c8e;
    ram_cell[     544] = 32'h02953623;
    ram_cell[     545] = 32'ha0e1c927;
    ram_cell[     546] = 32'hecc0fc76;
    ram_cell[     547] = 32'h3564beac;
    ram_cell[     548] = 32'h678ede98;
    ram_cell[     549] = 32'h56e97c95;
    ram_cell[     550] = 32'hf1d0314d;
    ram_cell[     551] = 32'h792b9480;
    ram_cell[     552] = 32'h1d20049e;
    ram_cell[     553] = 32'h9e699abe;
    ram_cell[     554] = 32'h28e9c11b;
    ram_cell[     555] = 32'hb2c23161;
    ram_cell[     556] = 32'hce5d476b;
    ram_cell[     557] = 32'hcafeb8df;
    ram_cell[     558] = 32'h780f8830;
    ram_cell[     559] = 32'ha72bb399;
    ram_cell[     560] = 32'h6583cc06;
    ram_cell[     561] = 32'hdcb4832e;
    ram_cell[     562] = 32'h1eb54e20;
    ram_cell[     563] = 32'h825d7e70;
    ram_cell[     564] = 32'h081a98a7;
    ram_cell[     565] = 32'h4d64feaf;
    ram_cell[     566] = 32'h6bac97db;
    ram_cell[     567] = 32'h315fe464;
    ram_cell[     568] = 32'h3db13dd7;
    ram_cell[     569] = 32'hbf75b5fa;
    ram_cell[     570] = 32'hc4fd71a0;
    ram_cell[     571] = 32'h4e46c4ee;
    ram_cell[     572] = 32'h6bf1d505;
    ram_cell[     573] = 32'hb851d757;
    ram_cell[     574] = 32'hcf51d39a;
    ram_cell[     575] = 32'h2ba4c653;
    ram_cell[     576] = 32'hcedb88da;
    ram_cell[     577] = 32'hcc5f94a3;
    ram_cell[     578] = 32'hf13fbc56;
    ram_cell[     579] = 32'hfe6b9b96;
    ram_cell[     580] = 32'h81142255;
    ram_cell[     581] = 32'hf2e15de4;
    ram_cell[     582] = 32'h67f68c38;
    ram_cell[     583] = 32'h385e7e72;
    ram_cell[     584] = 32'hf77e87dd;
    ram_cell[     585] = 32'h6e07fc04;
    ram_cell[     586] = 32'h3d9c95a0;
    ram_cell[     587] = 32'hb8641c65;
    ram_cell[     588] = 32'hda0d77d7;
    ram_cell[     589] = 32'hdb0671dc;
    ram_cell[     590] = 32'hff59ea80;
    ram_cell[     591] = 32'h3653d750;
    ram_cell[     592] = 32'h944464e3;
    ram_cell[     593] = 32'h348ef7d4;
    ram_cell[     594] = 32'hf4592db0;
    ram_cell[     595] = 32'h88ea0a0f;
    ram_cell[     596] = 32'h06e7a3d2;
    ram_cell[     597] = 32'h275b918f;
    ram_cell[     598] = 32'h245fced7;
    ram_cell[     599] = 32'he3dd304a;
    ram_cell[     600] = 32'hd8995e86;
    ram_cell[     601] = 32'h3220f0fb;
    ram_cell[     602] = 32'h06d4874a;
    ram_cell[     603] = 32'h50f9c137;
    ram_cell[     604] = 32'h5dd02c1a;
    ram_cell[     605] = 32'hbc9ab69c;
    ram_cell[     606] = 32'h464f4213;
    ram_cell[     607] = 32'heeafce53;
    ram_cell[     608] = 32'ha66e1673;
    ram_cell[     609] = 32'hc8d10312;
    ram_cell[     610] = 32'hc1d96fbc;
    ram_cell[     611] = 32'hba105722;
    ram_cell[     612] = 32'ha956f35e;
    ram_cell[     613] = 32'hb703d408;
    ram_cell[     614] = 32'h0cbdc5a1;
    ram_cell[     615] = 32'h4a5ba94b;
    ram_cell[     616] = 32'h69c02e39;
    ram_cell[     617] = 32'hccde6ab2;
    ram_cell[     618] = 32'hbb975665;
    ram_cell[     619] = 32'h1d9a6c64;
    ram_cell[     620] = 32'hcf415bd5;
    ram_cell[     621] = 32'hc8628108;
    ram_cell[     622] = 32'h87cf20c2;
    ram_cell[     623] = 32'hb4fcd40d;
    ram_cell[     624] = 32'hd97efd07;
    ram_cell[     625] = 32'h930cbb12;
    ram_cell[     626] = 32'hafb3f47e;
    ram_cell[     627] = 32'h8e541451;
    ram_cell[     628] = 32'h5ecb6db5;
    ram_cell[     629] = 32'h6f737804;
    ram_cell[     630] = 32'h1dae39b7;
    ram_cell[     631] = 32'hf17afc94;
    ram_cell[     632] = 32'h21c7e6c7;
    ram_cell[     633] = 32'h0e3d0640;
    ram_cell[     634] = 32'h7f892785;
    ram_cell[     635] = 32'h76cbd1bb;
    ram_cell[     636] = 32'hab9b1490;
    ram_cell[     637] = 32'h759a347a;
    ram_cell[     638] = 32'h8a1b8086;
    ram_cell[     639] = 32'h6dffb658;
    ram_cell[     640] = 32'h8295cbf4;
    ram_cell[     641] = 32'h5a70df7d;
    ram_cell[     642] = 32'h9810f270;
    ram_cell[     643] = 32'h2d2a318e;
    ram_cell[     644] = 32'hf6714113;
    ram_cell[     645] = 32'h31b18f60;
    ram_cell[     646] = 32'h76f3cd0e;
    ram_cell[     647] = 32'hf9833f8d;
    ram_cell[     648] = 32'hbcb67186;
    ram_cell[     649] = 32'hd331b35f;
    ram_cell[     650] = 32'h160820cf;
    ram_cell[     651] = 32'hc56868d6;
    ram_cell[     652] = 32'hc04c3b5e;
    ram_cell[     653] = 32'hc047c307;
    ram_cell[     654] = 32'h0e9300ec;
    ram_cell[     655] = 32'h7d3bf4b5;
    ram_cell[     656] = 32'h3af83868;
    ram_cell[     657] = 32'hf2554a7e;
    ram_cell[     658] = 32'h093f0a38;
    ram_cell[     659] = 32'h6cca0142;
    ram_cell[     660] = 32'h8bb13981;
    ram_cell[     661] = 32'h535fd199;
    ram_cell[     662] = 32'hb04e9840;
    ram_cell[     663] = 32'hbfa57a60;
    ram_cell[     664] = 32'h4514165b;
    ram_cell[     665] = 32'he4a12126;
    ram_cell[     666] = 32'hf3aa7e1d;
    ram_cell[     667] = 32'he7665b6d;
    ram_cell[     668] = 32'h87048194;
    ram_cell[     669] = 32'h54d003dc;
    ram_cell[     670] = 32'h21d40123;
    ram_cell[     671] = 32'h723c2b01;
    ram_cell[     672] = 32'hd85b6bf3;
    ram_cell[     673] = 32'hd7cf97e1;
    ram_cell[     674] = 32'h2236346a;
    ram_cell[     675] = 32'h652619dd;
    ram_cell[     676] = 32'hb9c69bfa;
    ram_cell[     677] = 32'h0cd655cf;
    ram_cell[     678] = 32'hc8904354;
    ram_cell[     679] = 32'h43b5026e;
    ram_cell[     680] = 32'h450105e6;
    ram_cell[     681] = 32'hfefc6b4f;
    ram_cell[     682] = 32'haa504987;
    ram_cell[     683] = 32'h9b20bbe4;
    ram_cell[     684] = 32'hccaceaa3;
    ram_cell[     685] = 32'h451bf978;
    ram_cell[     686] = 32'h493dd059;
    ram_cell[     687] = 32'hf41c0cd6;
    ram_cell[     688] = 32'hae277311;
    ram_cell[     689] = 32'h98dc1b9f;
    ram_cell[     690] = 32'h6b791b3c;
    ram_cell[     691] = 32'h1383da6c;
    ram_cell[     692] = 32'h03852af1;
    ram_cell[     693] = 32'hd40843ce;
    ram_cell[     694] = 32'hdadd3368;
    ram_cell[     695] = 32'he6758bde;
    ram_cell[     696] = 32'h56c0d9f0;
    ram_cell[     697] = 32'ha9887e41;
    ram_cell[     698] = 32'hc142157e;
    ram_cell[     699] = 32'h0f64289e;
    ram_cell[     700] = 32'hf2a86e84;
    ram_cell[     701] = 32'h03819d1e;
    ram_cell[     702] = 32'h3ac409e8;
    ram_cell[     703] = 32'h732d1ae2;
    ram_cell[     704] = 32'h5cb62280;
    ram_cell[     705] = 32'hc0d25e66;
    ram_cell[     706] = 32'h9b37d884;
    ram_cell[     707] = 32'h4ddaa36d;
    ram_cell[     708] = 32'h7c5d2a38;
    ram_cell[     709] = 32'h4ec5ddef;
    ram_cell[     710] = 32'h79d8076d;
    ram_cell[     711] = 32'hed1d05c9;
    ram_cell[     712] = 32'hb3568df9;
    ram_cell[     713] = 32'h27b0370b;
    ram_cell[     714] = 32'h851d3439;
    ram_cell[     715] = 32'h97b572d6;
    ram_cell[     716] = 32'ha6bf196f;
    ram_cell[     717] = 32'h62ebb962;
    ram_cell[     718] = 32'h62914ebf;
    ram_cell[     719] = 32'hb1dd253a;
    ram_cell[     720] = 32'h472ceab2;
    ram_cell[     721] = 32'h3d10f732;
    ram_cell[     722] = 32'h991de2e3;
    ram_cell[     723] = 32'hce67e066;
    ram_cell[     724] = 32'h8698db5b;
    ram_cell[     725] = 32'h42fe7b9b;
    ram_cell[     726] = 32'h4ff91606;
    ram_cell[     727] = 32'hb28d24d3;
    ram_cell[     728] = 32'h63a5fec3;
    ram_cell[     729] = 32'h1d67bd93;
    ram_cell[     730] = 32'h3b394827;
    ram_cell[     731] = 32'h77597b16;
    ram_cell[     732] = 32'h10fa6bff;
    ram_cell[     733] = 32'h26d287c4;
    ram_cell[     734] = 32'hfe6ac8b3;
    ram_cell[     735] = 32'hcbe73fe8;
    ram_cell[     736] = 32'h5c534d7b;
    ram_cell[     737] = 32'h29b57726;
    ram_cell[     738] = 32'he6c82b77;
    ram_cell[     739] = 32'h7e756296;
    ram_cell[     740] = 32'hcd22b2f6;
    ram_cell[     741] = 32'hca7f2569;
    ram_cell[     742] = 32'hefdd2159;
    ram_cell[     743] = 32'h3490194e;
    ram_cell[     744] = 32'h1886f26e;
    ram_cell[     745] = 32'h2c558a5c;
    ram_cell[     746] = 32'hd1e1d603;
    ram_cell[     747] = 32'h877260ba;
    ram_cell[     748] = 32'h7dbd0f22;
    ram_cell[     749] = 32'h01bdcc2c;
    ram_cell[     750] = 32'h9b617920;
    ram_cell[     751] = 32'hc6f27391;
    ram_cell[     752] = 32'hb22fa5bc;
    ram_cell[     753] = 32'ha0d6e48b;
    ram_cell[     754] = 32'hc37245b2;
    ram_cell[     755] = 32'h0e69edcd;
    ram_cell[     756] = 32'he2977084;
    ram_cell[     757] = 32'hadc666c6;
    ram_cell[     758] = 32'he888a0c5;
    ram_cell[     759] = 32'hc13f8f4d;
    ram_cell[     760] = 32'h0977d9f4;
    ram_cell[     761] = 32'h8c88c860;
    ram_cell[     762] = 32'h75bf818b;
    ram_cell[     763] = 32'h86584a7c;
    ram_cell[     764] = 32'h294a3d5f;
    ram_cell[     765] = 32'h41c69030;
    ram_cell[     766] = 32'h446a89fe;
    ram_cell[     767] = 32'h03e28378;
end

endmodule

